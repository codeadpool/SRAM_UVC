class sram_tx_monitor extends uvm_monitor;
  
endclass
