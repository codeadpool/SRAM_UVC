`include "sram_agent_pkg.sv"
package sram_seqs_pkg;
  import uvm_pkg::*;
  import sram_agent_pkg::*;
`include "sram_seq_lib.svh"
endpackage
