`include "sram_basic_test.sv"
`include "edge_seq_test.sv" 
`include "exhstve_seq_test.sv"
`include "rw_wr_test.sv"
