`include "sram_env_pkg.sv"
`include "uvm_macros.svh"
package sram_tests_pkg;
  import uvm_pkg::*;
  import sram_env_pkg::*;
  import sram_seqs_pkg::*;
  `include "sram_test_lib.svh"
endpackage
