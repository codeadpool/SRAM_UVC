package sram_package;
  parameter ADDR_WIDTH = 15;
  parameter DATA_WITDTH = 255;

endpackage
