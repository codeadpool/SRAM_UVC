`ifndef SRAM_DEFINES
`define SRAM_DEFINES
 `define ADDR_WIDTH 15
 `define NO_OF_TXS  20
`endif
